

module json2

pub type Map = map[string]Any
pub type Array = []Any

pub const (
	type_map = "map[string]json2.Any"
	type_array = "[]json2.Any"
)


